CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 70 2 150 10
176 80 1534 795
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 838 281 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.90056e-315 0
0
13 Logic Switch~
5 427 522 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3536 0 0
2
5.90056e-315 0
0
13 Logic Switch~
5 76 455 0 1 11
0 26
0
0 0 21344 0
1 7
-3 -16 4 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4597 0 0
2
5.90056e-315 0
0
13 Logic Switch~
5 69 264 0 1 11
0 27
0
0 0 21344 0
1 4
-3 -16 4 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3835 0 0
2
5.90056e-315 0
0
9 CA 7-Seg~
184 730 362 0 18 19
10 3 4 5 6 7 8 9 29 2
0 0 0 0 0 0 0 2 1
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3670 0 0
2
5.90056e-315 0
0
9 CA 7-Seg~
184 761 174 0 18 19
10 10 11 12 13 14 15 16 30 2
0 0 0 0 0 0 2 2 1
0
0 0 21104 0
7 AMBERCA
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5616 0 0
2
5.90056e-315 0
0
7 Pulser~
4 30 131 0 10 12
0 31 32 28 33 0 0 5 5 2
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
9323 0 0
2
5.90056e-315 0
0
6 74LS47
187 531 195 0 14 29
0 22 25 24 23 17 34 16 15 14
13 12 11 10 35
0
0 0 4832 0
6 74LS47
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
317 0 0
2
5.90056e-315 0
0
6 74LS47
187 537 380 0 14 29
0 21 20 19 18 17 36 9 8 7
6 5 4 3 37
0
0 0 4832 0
6 74LS47
-21 -60 21 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3108 0 0
2
5.90056e-315 0
0
6 74LS90
107 334 381 0 10 21
0 27 27 26 26 22 18 21 20 19
18
0
0 0 4832 0
6 74LS90
-21 -51 21 -43
2 U2
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
4299 0 0
2
5.90056e-315 0
0
6 74LS90
107 332 197 0 10 21
0 27 27 26 26 28 23 22 25 24
23
0
0 0 4832 0
6 74LS90
-21 -51 21 -43
2 U1
-7 -52 7 -44
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
9672 0 0
2
5.90056e-315 0
0
39
8 0 0 0 0 0 0 6 0 0 17 2
782 210
782 210
9 0 2 0 0 8192 0 5 0 0 3 4
730 326
730 292
859 292
859 281
9 1 2 0 0 8320 0 6 1 0 0 5
761 138
761 154
859 154
859 281
850 281
13 1 3 0 0 4224 0 9 5 0 0 5
575 398
675 398
675 437
709 437
709 398
12 2 4 0 0 4224 0 9 5 0 0 5
575 389
680 389
680 432
715 432
715 398
11 3 5 0 0 4224 0 9 5 0 0 5
575 380
685 380
685 427
721 427
721 398
10 4 6 0 0 4224 0 9 5 0 0 5
575 371
690 371
690 422
727 422
727 398
9 5 7 0 0 4224 0 9 5 0 0 5
575 362
695 362
695 417
733 417
733 398
8 6 8 0 0 4224 0 9 5 0 0 5
575 353
700 353
700 412
739 412
739 398
7 7 9 0 0 4224 0 9 5 0 0 5
575 344
705 344
705 407
745 407
745 398
13 1 10 0 0 4224 0 8 6 0 0 5
569 213
668 213
668 268
740 268
740 210
12 2 11 0 0 4224 0 8 6 0 0 5
569 204
673 204
673 263
746 263
746 210
11 3 12 0 0 4224 0 8 6 0 0 5
569 195
678 195
678 258
752 258
752 210
10 4 13 0 0 4224 0 8 6 0 0 5
569 186
683 186
683 253
758 253
758 210
9 5 14 0 0 4224 0 8 6 0 0 5
569 177
688 177
688 248
764 248
764 210
8 6 15 0 0 4224 0 8 6 0 0 5
569 168
693 168
693 243
770 243
770 210
7 7 16 0 0 4240 0 8 6 0 0 6
569 159
698 159
698 238
782 238
782 210
776 210
5 0 17 0 0 4096 0 9 0 0 19 2
505 416
448 416
5 1 17 0 0 8320 0 8 2 0 0 4
499 231
448 231
448 522
439 522
10 4 18 0 0 4224 0 10 9 0 0 4
366 408
476 408
476 371
505 371
9 3 19 0 0 4224 0 10 9 0 0 4
366 390
486 390
486 362
505 362
8 2 20 0 0 4224 0 10 9 0 0 4
366 372
481 372
481 353
505 353
7 1 21 0 0 4224 0 10 9 0 0 4
366 354
486 354
486 344
505 344
5 0 22 0 0 8320 0 10 0 0 28 5
296 399
294 399
294 150
399 150
399 170
10 4 23 0 0 4224 0 11 8 0 0 4
364 224
481 224
481 186
499 186
9 3 24 0 0 4224 0 11 8 0 0 4
364 206
491 206
491 177
499 177
8 2 25 0 0 4224 0 11 8 0 0 4
364 188
486 188
486 168
499 168
7 1 22 0 0 0 0 11 8 0 0 4
364 170
491 170
491 159
499 159
6 10 18 0 0 0 0 10 10 0 0 6
296 408
292 408
292 423
374 423
374 408
366 408
6 10 23 0 0 0 0 11 11 0 0 6
294 224
290 224
290 239
372 239
372 224
364 224
4 0 26 0 0 4096 0 10 0 0 32 3
302 381
201 381
201 372
3 0 26 0 0 4096 0 10 0 0 34 3
302 372
98 372
98 455
4 0 26 0 0 0 0 11 0 0 34 3
300 197
187 197
187 188
3 1 26 0 0 8320 0 11 3 0 0 4
300 188
102 188
102 455
88 455
2 0 27 0 0 4096 0 11 0 0 36 3
300 179
189 179
189 170
1 0 27 0 0 4096 0 11 0 0 38 4
300 170
95 170
95 264
90 264
2 0 27 0 0 0 0 10 0 0 38 3
302 363
205 363
205 354
1 1 27 0 0 4224 0 10 4 0 0 4
302 354
90 354
90 264
81 264
3 5 28 0 0 4224 0 7 11 0 0 4
54 122
286 122
286 215
294 215
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
